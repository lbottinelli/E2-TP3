// Define Key Code Constants

parameter KEY_1 = 4'b 0000;
parameter KEY_2 = 4'b 0001;
parameter KEY_3 = 4'b 0010;
parameter KEY_A = 4'b 0011;
parameter KEY_4 = 4'b 0100;
parameter KEY_5 = 4'b 0101;
parameter KEY_6 = 4'b 0110;
parameter KEY_B = 4'b 0111;
parameter KEY_7 = 4'b 1000;
parameter KEY_8 = 4'b 1001;
parameter KEY_9 = 4'b 1010;
parameter KEY_C = 4'b 1011;
parameter KEY_ASS = 4'b 1100;
parameter KEY_0 = 4'b 1101;
parameter KEY_HASH = 4'b 1110;
parameter KEY_D = 4'b 1111;
