module fsm_module (clk, enable_in, reset_in, out);
    input wire clk, enable_in, reset_in;
    output wire [3:0] out;

    always @(posedge clk) begin
        
    end

endmodule